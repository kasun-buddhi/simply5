////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
// Author       : kasun buddhi
// email        : kasun@kasunbuddhi.com
// date         : 2024.07.15
// file         : core.sv
// Description  : this is the core which instantiate all other components of the core here 
//                ex : alu, control units, decoder, accumilator 
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////

module core (

);

endmodule : core