////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
// Author       : kasun buddhi
// email        : kasun@kasunbuddhi.com
// date         : 2024.07.18
// file         : decoder.sv
// Description  : this is the decoder
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////